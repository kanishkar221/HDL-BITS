module top_module( 
    input a,b,c,
    output w,x,y,z );
    
    assign w = a;
	  assign y = b;
   	assign x = b;
    assign z = c;
endmodule
