module top_module(
    input clk,
    input in,
    input reset,    // Synchronous reset
    output done
);
    parameter IDLE = 3'b000;
	  parameter START = 3'b001;
	  parameter RECEIVE = 3'b010;
	  parameter WAIT = 3'b011;
	  parameter STOP = 3'b100;

	  reg [2:0] state, next;
	  reg [3:0] i;

	  always @(*) begin
		  case(state)
			  IDLE  : next = (in) ? IDLE : START;
			  START : next = RECEIVE;
			  RECEIVE : begin
				  if (i == 8) begin
					  if (in) next = STOP;
					  else next = WAIT;
				  end 
				  else next = RECEIVE;			
			  end
			  WAIT : next = (in) ? IDLE : WAIT;
			  STOP : next = (in) ? IDLE : START;
		  endcase
	  end

	  always @(posedge clk) begin
		  if(reset) state <= IDLE;
		  else state <= next;
	  end

	  always @(posedge clk) begin
		  if (reset) begin
			  done <= 0;
			  i <= 0;
		  end
		  else begin
			  case(next) 
				  RECEIVE : begin
					  done <= 0;
					  i = i + 1;
				  end
				  STOP : begin
					  done <= 1;
					  i <= 0;
				  end
				  default : begin
					  done <= 0;
					  i <= 0;
				  end
			  endcase
		  end
	  end
endmodule
