module top_module(
    output zero
);// Module body
    assign zero = 1'b0;

endmodule

